library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity mine2 is
  generic(ID: integer := 0);
  port(
    reset: in std_logic; 
    clk: in std_logic; -- 50 MHz clock; used for count-down timers only
    countdown_timer_tick: in std_logic; -- used by 2 sec and 4 sec countdown timers
    TIME_TICK: in std_logic; -- clock of 30 cycles per second
    x0, y0: in std_logic_vector(9 downto 0); -- location where mine is planted
    MINE2_PLANT: in std_logic;
    MINE2_RECYCLE: in std_logic;
    MINE2_IMG: out std_logic; -- event generated to Tunnel    
    mine2_bmp_overlaps_ship_bmp: in std_logic; -- from checker of collision with ship, from Tunnel
    HIT_MINE2: out std_logic; -- event generated to Ship
    mine2_bmp_overlaps_missile_bmp: in std_logic; -- from checker of collision with missile
    mine2_hit_1st_time: out std_logic; -- event generated by mine2 for missile, passed via Tunnel
    DESTROYED_MINE2: out std_logic; -- event generated to Missile
    EXPLOSION_MINE2: out std_logic; -- event generated to Tunnel
    exit_action: in std_logic; -- from Player
    MINE2_DISABLED: out std_logic; -- event generated to Tunnel
    mine2_id: out std_logic_vector(2 downto 0); -- info passed with event MINE2_DISABLED
    x, y: out std_logic_vector(9 downto 0); -- coordinates passed with events posted
    mine2_explosion_size: out std_logic_vector(9 downto 0) -- passed with event EXPLOSION_MINE2
  );
end mine2;


architecture UML_ARCHITECTURE of mine2 is

  type SUPERSTATE_TYPE_MINE2 is (USED, UNUSED);
  type STATE_TYPE_MINE2 is (Planted, Exploding);
  signal superstate_reg, superstate_next: SUPERSTATE_TYPE_MINE2;
  signal state_reg, state_next: STATE_TYPE_MINE2;
  -- coordinates where mine is planted;
  signal x_reg, x_next: unsigned(9 downto 0);
  signal y_reg, y_next: unsigned(9 downto 0);
  signal local_ctr_reg, local_ctr_next: unsigned(7 downto 0); -- local counter; count TIME_TICK 30 times (i.e., 1 sec) and increment score
  signal exp_ctr_reg, exp_ctr_next: unsigned(9 downto 0); -- explosion counter 
  signal missile_hits_ctr_reg, missile_hits_ctr_next: unsigned(1 downto 0); -- when mine is hit twice only it explodes  

  constant MAX_X: integer:=640;
  constant MAX_Y: integer:=480;
  constant MINE2_HEIGHT: integer:=32;
  constant MINE2_DELTA_V: integer:=1; 
  signal timer_2sec_start, timer_2sec_up: std_logic;
  
  
  begin
    
    -- state register; process #1
    process (TIME_TICK, reset)
    begin
      if (reset = '1') then 
        superstate_reg <= UNUSED;
        state_reg <= Planted;
        --x_reg <= to_unsigned(MAX_X,10); -- place mine20 in the middle of screen on x axis;
        --y_reg <= to_unsigned((MAX_Y-MINE2_HEIGHT)/2,10); -- place mine20 in the middle of screen on y axis;
        x_reg <= unsigned(x0);
        y_reg <= unsigned(y0);
        local_ctr_reg <= (OTHERS=>'0');
        exp_ctr_reg <= (OTHERS=>'0');
        missile_hits_ctr_reg <= "00";
      elsif (TIME_TICK' event and TIME_TICK = '1') then 
        superstate_reg <= superstate_next;
        state_reg <= state_next;
        x_reg <= x_next;
        y_reg <= y_next;
        exp_ctr_reg <= exp_ctr_next;
        local_ctr_reg <= local_ctr_next;
        missile_hits_ctr_reg <= missile_hits_ctr_next;
      end if;
    end process;    
    
    
    -- next state and output logic; process #2
    process (superstate_reg, state_reg, MINE2_PLANT, MINE2_RECYCLE, 
      mine2_bmp_overlaps_ship_bmp, mine2_bmp_overlaps_missile_bmp, 
      exit_action)
    begin
      -- default initializations
      superstate_next <= superstate_reg;
      state_next <= state_reg;
      x_next <= x_reg;
      y_next <= y_reg;
      exp_ctr_next <= exp_ctr_reg;
      local_ctr_next <= local_ctr_reg;
      missile_hits_ctr_next <= missile_hits_ctr_reg;
      mine2_hit_1st_time <= '0';
      MINE2_IMG <= '0';
      HIT_MINE2 <= '0';
      DESTROYED_MINE2 <= '0';
      EXPLOSION_MINE2 <= '0';
      MINE2_DISABLED <= '0';
      timer_2sec_start <='0';      
  
      case superstate_reg is 
        --=====================================================================
        when UNUSED => -- superstate
          if MINE2_PLANT = '1' then
            superstate_next <= USED;
            state_next <= Planted;
            x_next <= unsigned(x0);
            y_next <= unsigned(y0);
            missile_hits_ctr_next <= "00"; --reset hits counter, in case it was incremented once only and then got out of screen
          end if;  
        --=====================================================================
        when USED => -- superstate; 
          if exit_action = '1' then 
            MINE2_DISABLED <= '1'; -- tell the Tunnel object
            superstate_next <= UNUSED;
          end if;
          if MINE2_RECYCLE = '1' then
            superstate_next <= UNUSED;
          end if;
          -- [case statement] for the inner states of "USED" superstate
          case state_reg is 
            --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
            when Planted =>
              MINE2_IMG <= '1';
              if (x_reg >= MINE2_DELTA_V) then -- I can continue to move to the left a "delta v" on screen          
                x_next <= x_reg - MINE2_DELTA_V; -- moving to the left with Tunnel creates the illusion of Ship moving to right
              else -- if I subtractd MINE2_DELTA_V pixels I would place left edge of mine outside screen on left; I work with unsigned!
                superstate_next <= UNUSED; -- mine out of boundary of screen
              end if;          
              if (mine2_bmp_overlaps_missile_bmp = '1') then 
                if (missile_hits_ctr_reg=1) then -- this is alread the 2nd hit by a missile; done, explode
                  DESTROYED_MINE2 <= '1'; -- generate event to Missile
                  state_next <= Exploding; 
                  exp_ctr_next <= (OTHERS=>'0'); -- clear explosion counter
                  timer_2sec_start <='1'; -- start cowntdown counter 2 sec
                  missile_hits_ctr_next <= "00"; --reset hits counter
                else 
                  missile_hits_ctr_next <= missile_hits_ctr_reg + 1; -- increment hits counter
                  mine2_hit_1st_time <= '1';
                end if;
              end if;
              if (mine2_bmp_overlaps_ship_bmp = '1') then 
                HIT_MINE2 <= '1'; -- generate event to Ship
                superstate_next <= UNUSED; 
              end if;            
            --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~                
            when Exploding =>
              EXPLOSION_MINE2 <= '1'; -- post event to Tunnel
              -- wait for 2 sec to display exploding ship
              if timer_2sec_up='1' then
                superstate_next <= UNUSED; 
              end if;               
            --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
          end case;     
        --=====================================================================  
      end case;
    end process;
 
  -- coordinates passed with events 
  x <= std_logic_vector(x_reg);
  y <= std_logic_vector(y_reg); 
    
  mine2_id <= std_logic_vector(to_unsigned(ID,3));
  
  -- instantiate countdown timer
  timer_2sec_mine2_U0: entity work.timer
    generic map(W=>6) -- 2 seconds timer
    port map(clk=>clk, reset=>reset,
            timer_tick=>countdown_timer_tick,
            timer_start=>timer_2sec_start,
            timer_up=>timer_2sec_up);
            
end UML_ARCHITECTURE;  
