library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity tunnel_and_graph is
   port(
      clk, clk_10Hz: in std_logic; -- clk is 50 MHz 
      countdown_timer_tick: in std_logic; -- used by 2 sec and 4 sec countdown timers
      pixel_tick: in std_logic; -- comes from vga_sync entity from top level
      reset: in std_logic;     
      in_state_new_game: out std_logic; -- is Tunnel in state NEW_GAME?
      in_state_game_over_message: out std_logic; -- is Tunnel in state GAME_OVER_MESSAGE?
      vsync: in std_logic; -- will be used as 1/30 sec TIME_TICK
      btn: std_logic_vector(2 downto 0); -- KEY2: fire Missile; KEY1,0: Ship down/up;
      pixel_x,pixel_y: in std_logic_vector(9 downto 0);
      graph_on: out std_logic;
      score: out std_logic_vector(19 downto 0); -- will be passed to game_text entity at top level
      rgb: out std_logic_vector(2 downto 0) -- this is graphics rgb signal; will be muxed with text rgb at top level
   );
end tunnel_and_graph;


architecture arch of tunnel_and_graph is
  constant MAX_X: integer:=640;
  constant MAX_Y: integer:=480;
  constant SCORE_DELTA_FOR_MINE1: integer:=20;
  constant SCORE_DELTA_FOR_MINE2: integer:=50;
  
  constant NO_MINE1_PLANT_ZONE_XL: integer:=100;
  constant NO_MINE1_PLANT_ZONE_XR: integer:=440;
  constant NO_MINE2_PLANT_ZONE_XL: integer:=300;
  constant NO_MINE2_PLANT_ZONE_XR: integer:=640;
  
  signal pix_x, pix_y: unsigned(9 downto 0);

  signal timer_4sec_start, timer_4sec_up: std_logic;
  signal game_exit_from_user: std_logic; -- from Player
  
  signal tunnel_rgb: std_logic_vector(2 downto 0);
  signal ship_rgb, ship_expl_rgb: std_logic_vector(2 downto 0);
  signal missile_rgb, missile_expl_rgb: std_logic_vector(2 downto 0);
  signal mine10_rgb, mine10_expl_rgb: std_logic_vector(2 downto 0);
  signal mine20_rgb, mine20_expl_rgb: std_logic_vector(2 downto 0);
  
 
  -- MINES
  constant MINE1_WIDTH: integer:=24; -- mine type 1
  constant MINE1_HEIGHT: integer:=24;
  constant MINE2_WIDTH: integer:=32; -- mine type 2
  constant MINE2_HEIGHT: integer:=32;
  
  signal seed_for_LFSR: unsigned(9 downto 0);   
  signal x_rand_lfsr_mine10, y_rand_lfsr_mine10: unsigned(9 downto 0); -- random numbers generated by LFSRs
  signal x_rand_lfsr_mine20, y_rand_lfsr_mine20: unsigned(9 downto 0); -- random numbers generated by LFSRs
  signal mine10_x_rand_reg, mine10_y_rand_reg: unsigned(9 downto 0); -- random numbers that qualify for planting mine10
  signal mine10_x_rand_next, mine10_y_rand_next: unsigned(9 downto 0);
  signal mine20_x_rand_reg, mine20_y_rand_reg: unsigned(9 downto 0); -- random numbers that qualify for planting mine20
  signal mine20_x_rand_next, mine20_y_rand_next: unsigned(9 downto 0);
  
	type STATE_TYPE_PLANTING_MINES is (PLANT_PAUSE, PLANT_MINE1, PLANT_MINE2);
  signal plant_mine_state_reg, plant_mine_state_next: STATE_TYPE_PLANTING_MINES;
  
  
  -- mine1
  signal mine10_x_l, mine10_x_r: unsigned(9 downto 0);
  signal mine10_y_t, mine10_y_b: unsigned(9 downto 0);
  signal mine10_x_rand, mine10_y_rand: unsigned(9 downto 0); -- location where mine is planted randomly eventually  
  signal mine10_x_reg, mine10_x_next: unsigned(9 downto 0); -- location of mine on screen for display purposes 
  signal mine10_y_reg, mine10_y_next: unsigned(9 downto 0); 
  signal bbox_mine10_on, actual_mine10_on: std_logic; 
  signal bbox_expanded_mine10_on: std_logic; -- area to avoid to place the other mine;
  signal mine10_curr_x: std_logic_vector(9 downto 0); -- coordinates passed with events posted
  signal mine10_curr_y: std_logic_vector(9 downto 0); -- coordinates passed with events posted 
  signal plant_mine10: std_logic;
  signal recycle_mine10: std_logic;
  signal mine10_is_planted: std_logic; -- event generated to Tunnel  
  signal ship_hit_mine10_ev, ship_hit_mine10_ev_recorded: std_logic; -- event generated to Ship
  signal ship_hit_mine_from_mine10: std_logic; -- from mines to ship
  signal missile_hit_mine10_ev, missile_hit_mine10_ev_recorded: std_logic; -- from checker of collision with missile 
  signal missile_destroyed_mine10: std_logic; -- event generated to Missile
  signal explode_mine10: std_logic; -- event generated to Tunnel  
  signal mine10_disabled: std_logic; -- event generated to Tunnel
  signal mine10_id: std_logic_vector(2 downto 0); -- info passed with event MINE1_DISABLED
  signal mine10_explosion_size : std_logic_vector(9 downto 0); -- passed with event EXPLOSION_MINE1

  
  -- mine2
  signal mine20_x_l, mine20_x_r: unsigned(9 downto 0);
  signal mine20_y_t, mine20_y_b: unsigned(9 downto 0);
  signal mine20_x_rand, mine20_y_rand: unsigned(9 downto 0); -- location where mine is planted randomly eventually  
  signal mine20_x_reg, mine20_x_next: unsigned(9 downto 0); -- location of mine on screen for display purposes 
  signal mine20_y_reg, mine20_y_next: unsigned(9 downto 0); 
  signal bbox_mine20_on, actual_mine20_on: std_logic; 
  signal bbox_expanded_mine20_on: std_logic; -- area to avoid to place the other mine;
  signal mine20_curr_x: std_logic_vector(9 downto 0); -- coordinates passed with events posted
  signal mine20_curr_y: std_logic_vector(9 downto 0); -- coordinates passed with events posted 
  signal plant_mine20: std_logic;
  signal recycle_mine20: std_logic;
  signal mine20_is_planted: std_logic; -- event generated to Tunnel  
  signal ship_hit_mine20_ev, ship_hit_mine20_ev_recorded: std_logic; -- event generated to Ship
  signal ship_hit_mine_from_mine20: std_logic; -- from mines to ship
  signal missile_hit_mine20_ev, missile_hit_mine20_ev_recorded: std_logic; -- from checker of collision with missile 
  signal missile_destroyed_mine20: std_logic; -- event generated to Missile
  signal explode_mine20: std_logic; -- event generated to Tunnel
  signal missile_hit_mine20_1st_time: std_logic; -- event generated by mine20 for missile via Tunnel
  signal mine20_disabled: std_logic; -- event generated to Tunnel
  signal mine20_id: std_logic_vector(2 downto 0); -- info passed with event MINE2_DISABLED
  signal mine20_explosion_size : std_logic_vector(9 downto 0); -- passed with event EXPLOSION_MINE2
  
  -- mine 1
  type MINE1_ROM_TYPE is array (0 to 23) of std_logic_vector(23 downto 0);
  constant mine10_bmp: MINE1_ROM_TYPE :=
  (
    "000000000000011000000000", --0
    "000000111000111100000000", --1
    "000001111000111100000000", --2
    "000001111111111100000000", --3
    "000001111111111111001100", --4
    "000001111111111111111110", --5
    "000011111111111111111110", --6
    "001111100011111111111110", --7
    "111111000001111111111000", --8
    "111111000001111111111000", --9
    "111111100011111111111100", --10
    "011111111111111111111100", --11
    "001111111111111111111100", --12
    "001111111111111111111111", --13
    "001111111111111111111111", --14
    "001111111111111111111111", --15
    "011111111111111111111000", --16
    "011111111111111111110000", --17
    "011111111111111111110000", --18
    "001101111111111111100000", --19
    "000000111111111111110000", --20
    "000000001111111011110000", --21
    "000000001110000011100000", --22
    "000000001110000000000000"  --23
  );
  signal mine10_rom_addr: unsigned(4 downto 0);
  signal mine10_rom_col: unsigned(4 downto 0);
  signal mine10_rom_data: std_logic_vector(23 downto 0);
  signal mine10_rom_bit: std_logic;

  -- mine 2
  type MINE2_ROM_TYPE is array (0 to 31) of std_logic_vector(31 downto 0);
  constant mine20_bmp: MINE2_ROM_TYPE :=
  (
    "00000000000110000001100000000000", --0
    "00000000011100000000111000000000", --1
    "00000000111000000000011000000000", --2
    "00000000110000000000011100000000", --3
    "00000001110000000000001110000000", --4
    "00000001110011111110001110000000", --5
    "00000001110111111111101110000000", --6
    "00000011111111111111111110000000", --7
    "00000011111111111111111110000000", --8
    "00000011111111111111111110000000", --9
    "00000001111111111111111110000000", --10
    "00000011111111111111111111000000", --11
    "00001111111111111111111111110000", --12
    "00011111111111111111111111111100", --13
    "00111111100111111111001111111110", --14
    "01111111100011111110001111111110", --15
    "01111000111101111101111100001111", --16
    "11100000011111111111111100000111", --17
    "11000000011111011011111100000011", --18
    "11000000011111111111111100000001", --19
    "10000000001101111111011000000001", --20
    "10000000000001011101000000000001", --21
    "10000000000001011101000000000001", --22
    "00000000000001011101000000000000", --23
    "00000000000001011101000000000000", --24
    "00000000000001011101000000000000", --25
    "00000000000001011101000000000000", --26
    "00000000000011111111100000000000", --27
    "00000000000111111111110000000000", --28
    "00000000001111111111111000000000", --29
    "00111111111111100011111111111100", --30
    "00001111111110000000111111110000"  --31
  );
  signal mine20_rom_addr: unsigned(4 downto 0);
  signal mine20_rom_col: unsigned(4 downto 0);
  signal mine20_rom_data: std_logic_vector(31 downto 0);
  signal mine20_rom_bit: std_logic;
  

  -- Missile related signals
  constant MISSILE_WIDTH: integer:=16; 
  constant MISSILE_HEIGHT: integer:=8; 
  signal missile_x_l, missile_x_r: unsigned(9 downto 0);
  signal missile_y_t, missile_y_b: unsigned(9 downto 0);
  signal missile_x_reg, missile_x_next: unsigned(9 downto 0);
  signal missile_y_reg, missile_y_next: unsigned(9 downto 0);
  signal bbox_missile_on, actual_missile_on: std_logic; 
  constant MISSILE_VELOCITY: unsigned(9 downto 0) :=to_unsigned(2,10); 
  signal missile_curr_x: std_logic_vector(9 downto 0); -- coordinates passed with events posted by missile 
  signal missile_curr_y: std_logic_vector(9 downto 0);
  signal missile_hit_mine : std_logic; -- event posted by Tunnel 
  signal missile_destroyed_mine: std_logic; -- event posted by Tunnel 
  signal missile_hit_wall_ev : std_logic; -- event posted by Tunnel  
  signal missile_IMG_ev : std_logic; -- event posted to Tunnel
  signal score_delta_val_from_missile: std_logic_vector(19 downto 0);
  signal explode_missile: std_logic; -- event posted to Tunnel
  signal missile_explosion_size: std_logic_vector(9 downto 0); -- passed with event EXPLOSION_MISSILE 
  signal missile_is_flying: std_logic;
  
  type MISSILE_ROM_TYPE is array (0 to 7) of std_logic_vector(15 downto 0);
  constant missile_bmp: MISSILE_ROM_TYPE :=
  (
    "1111111111111000",
    "1111111111111100",
    "1111111111111110",
    "1111111111111111", 
    "1111111111111111",
    "1111111111111110",
    "1111111111111100",
    "1111111111111000"
  );
  signal missile_rom_addr: unsigned(2 downto 0);
  signal missile_rom_col: unsigned(3 downto 0);
  signal missile_rom_data: std_logic_vector(15 downto 0);
  signal missile_rom_bit: std_logic;


  -- Ship related signals
  constant SHIP_WIDTH : integer:=48;
  constant SHIP_HEIGHT : integer:=32;
  constant SHIP_DELTA_V: integer:=2;
  signal TIME_TICK: std_logic; -- tick at which the Ship moves, ship tick
  signal ship_x_l, ship_x_r : unsigned(9 downto 0);
  signal ship_y_t, ship_y_b : unsigned(9 downto 0);
  signal ship_x_reg, ship_x_next: unsigned(9 downto 0);
  signal ship_y_reg, ship_y_next: unsigned(9 downto 0);
  signal bbox_ship_on, actual_ship_on: std_logic;
  
  signal player_fire_missile: std_logic;
  signal player_ship_move: std_logic; -- event that comes with coordinates info
  signal take_off_ev : std_logic; -- event generated by Tunnel when Player starts game
  signal score_total_val : std_logic_vector(19 downto 0); -- ship total accumulated score value, passed with event SCORE 
  signal score_ev : std_logic; -- event generated
  signal ship_curr_x : std_logic_vector(9 downto 0); -- passed with event SHIP_IMG
  signal ship_curr_y : std_logic_vector(9 downto 0); -- passed with event SHIP_IMG
  signal ship_IMG_ev : std_logic; -- event posted to Tunnel
  signal ship_hit_mine : std_logic; -- event posted by Tunnel; either mine1 OR mine2; ship explodes anyways
  signal mine_type_hit : std_logic_vector(1 downto 0); -- actually we have just 2 types of mines
  signal ship_hit_wall_ev : std_logic; -- event posted by Tunnel
  signal fire_missile : std_logic; -- event posted to Missile; includes x,y too
  signal destroyed_mine_ev : std_logic; -- event from Missile to Ship
  signal score_delta_destroyed_mine_1_or_2 : std_logic_vector(19 downto 0); -- how much to add to local score when mine is destroyed
  signal explode_ship: std_logic; -- event posted to Tunnel
  signal ship_explosion_size : std_logic_vector(9 downto 0); -- passed with event EXPLOSION_SHIP
  signal game_over_from_ship: std_logic;
  signal ship_is_flying: std_logic;
  
  -- ROM Type for Ship
  type SHIP_ROM_TYPE is array (0 to 31) of std_logic_vector (47 downto 0);
  constant ship_bmp: SHIP_ROM_TYPE := 
    (
    "000000000000111111000011111100000000000000000000", --0
    "000000000111111111111111111111000000000000000000", --1
    "000000011111111111111111111111111000000000000000", --2
    "000000111111111111111111111111111111000000000000", --3
    "000001111111111111111111111111111111111000000000", --4
    "000011111111111111111111111111111111111111000000", --5
    "000111111111111111111111111111111111111111111000", --6
    "001111111111111111111111111111111111111111111111", --7
    "011111111111111111111111111111111111111111111111", --8
    "011111111111111111111111111111111111111111111111", --9
    "011111111111111100000001111111111111111111111111", --10
    "111111111111111000111000011111111111111111111111", --11
    "111111111111110011111110000000000000000000000000", --12
    "111111111111100111111111000111111111111100000000", --13
    "111111111111100111111111100111111111111100000000", --14
    "111111111111000111111111100111111111111100000000", --15
    "111111111111100111111111100111111111111100000000", --16
    "111111111111100111111111000111111111111100000000", --17
    "111111111111110011111111000111111111111100000000", --18
    "111111111111111000111100000000000000000000000000", --19
    "111111111111111100000000111111111111111111111111", --20
    "011111111111111111111111111111111111111111111111", --21
    "011111111111111111111111111111111111111111111111", --22
    "001111111111111111111111111111111111111111111111", --23
    "000111111111111111111111111111111111111111111111", --24
    "000011111111111111111111111111111111111111111000", --25
    "000001111111111111111111111111111111111100000000", --26
    "000000111111111111111111111111110000000000000000", --27
    "000000011111111111111111111111111111111100000000", --28
    "000000000111111111111111111111111111111100000000", --29
    "000000000001111111000001111111111111111100000000", --30
    "000000000000000000000000000001111111111100000000"  --31
    );
  signal ship_rom_addr: unsigned(4 downto 0);
  signal ship_rom_col: unsigned(5 downto 0);
  signal ship_rom_data: std_logic_vector(47 downto 0);
  signal ship_rom_bit: std_logic;  
  
  
  -- EXPLOSIONS signals
  constant MISSILE_EXPL_WIDTH: integer:=32; 
  constant MISSILE_EXPL_HEIGHT: integer:=24; 
  -- missile - explosion is with larger bbox than missile itself, so I need to keep track of these:
  signal missile_expl_x_l, missile_expl_x_r: unsigned(9 downto 0);
  signal missile_expl_y_t, missile_expl_y_b: unsigned(9 downto 0);
  --location of impact with wall; "frozen" on Tunnel
  --so that missile explosion stays at place of collision and
  --does not continue to move to the right
  signal missile_x0_explosion_reg, missile_x0_explosion_next: unsigned(9 downto 0); 
  signal bbox_missile_expl_on, actual_missile_expl_on: std_logic; 
  signal missile_hit_wall_ev_recorded: std_logic;
  --ship
  signal ship_x0_explosion_reg, ship_x0_explosion_next: unsigned(9 downto 0); 
  signal actual_ship_expl_on: std_logic;
  signal ship_hit_wall_ev_recorded: std_logic; 
  --mine10
  signal mine10_expl_x_l, mine10_expl_x_r: unsigned(9 downto 0);
  signal mine10_expl_y_t, mine10_expl_y_b: unsigned(9 downto 0);
  signal bbox_expl_mine10_on, actual_mine10_expl_on: std_logic; 
  signal mine10_x0_explosion_reg, mine10_x0_explosion_next: unsigned(9 downto 0);   
  --mine20
  signal mine20_expl_x_l, mine20_expl_x_r: unsigned(9 downto 0);
  signal mine20_expl_y_t, mine20_expl_y_b: unsigned(9 downto 0);
  signal bbox_expl_mine20_on, actual_mine20_expl_on: std_logic; 
  signal mine20_x0_explosion_reg, mine20_x0_explosion_next: unsigned(9 downto 0); 
  
  -- ROM Type for Ship EXPLOSION
  type SHIP_EXPLOSION_ROM_TYPE is array (0 to 31) of std_logic_vector (47 downto 0);
  constant ship_expl_bmp: SHIP_EXPLOSION_ROM_TYPE := 
    (       
    "000000000000000000000000000000011000000000000000", --0
    "000000000000000000000000000000111000000000000000", --1
    "000000000000000000000000000001111000000000000000", --2
    "011000000000000000110000000011111000000000000000", --3
    "011111000000000000111000000111111000000000000000", --4
    "000111110000000001111100000111111000000000000000", --5
    "000011111110000001111110001111110000000111000000", --6
    "000001111111100001111111011111111111111110000000", --7
    "000000111111111111111111111111111111111100000000", --8
    "000000011111111111111111111111111111111100000000", --9
    "000000001111111111111111111111111111111000000000", --10
    "000000011111111111111111111111111111111111111100", --11
    "111111111111111111111111111111111111111111111110", --12
    "111111111111111111111111111111111111111111111100", --13
    "001111111111111111111111111111111111111111110000", --14
    "000011111111111111111111111111111111111110000000", --15
    "000001111111111111111111111111111111111111100000", --16
    "000000011111111111111111111111111111111111111000", --17
    "000000111111111111111111111111111111111111111110", --18
    "000011111111111111111111111111111111111111111111", --19
    "001111111111111111111111111111111111111000000000", --20
    "111111111111111111111111111111111111111000000000", --21
    "000000000000111111111111111111111111111100000000", --22
    "000000000001111111111111111111110111111100000000", --23
    "000000000001111111111110011111100001111100000000", --24
    "000000000001110001111110001111100000011110000000", --25
    "000000000001000000111110001111100000001110000000", --26
    "000000000000000000111100000111100000000000000000", --27
    "000000000000000000111100000011100000000000000000", --28
    "000000000000000000111000000001000000000000000000", --29
    "000000000000000000111000000000000000000000000000", --30
    "000000000000000000110000000000000000000000000000"  --31
    );
  signal ship_expl_rom_addr: unsigned(4 downto 0);
  signal ship_expl_rom_col: unsigned(5 downto 0);
  signal ship_expl_rom_data: std_logic_vector(47 downto 0);
  signal ship_expl_rom_bit: std_logic;   
  
  -- ROM Type for Missile EXPLOSION (when it hits the walls)
  type MISSILE_EXPLOSION_ROM_TYPE is array (0 to 23) of std_logic_vector (31 downto 0);
  constant missile_expl_bmp: MISSILE_EXPLOSION_ROM_TYPE := 
    (       
    "00000000000000000000001000000000", --0
    "00000000000000000000011000000000", --1
    "00000000000010000000111000000000", --2
    "11000000000111000001111000000000", --3
    "11111000000111100011111000000000", --4
    "01111110000111110111111111111100", --5
    "00111111111111111111111111111000", --6
    "00011111111111111111111111110000", --7
    "00001111111111111111111111111111", --8
    "11111111111111111111111111111111", --9
    "11111111111111111111111111111111", --10
    "00111111111111111111111111111100", --11
    "00011111111111111111111111111000", --12
    "00011111111111111111111111111111", --13
    "01111111111111111111111111111110", --14
    "11111111111111111111111111110000", --15
    "11110001111111111111111111110000", --16
    "00000011111111111111110111111000", --17
    "00000011111111110111110001111000", --18
    "00000011000111100011110000111100", --19
    "00000000000111100011110000001100", --20
    "00000000000111000001100000000000", --21
    "00000000000011000000100000000000", --22
    "00000000000011000000000000000000"  --23
    );
  signal missile_expl_rom_addr: unsigned(4 downto 0);
  signal missile_expl_rom_col: unsigned(4 downto 0);
  signal missile_expl_rom_data: std_logic_vector(31 downto 0);
  signal missile_expl_rom_bit: std_logic;  
  
  -- mine1 explosion
  type MINE1_EXPL_ROM_TYPE is array (0 to 23) of std_logic_vector(23 downto 0);
  constant mine10_expl_bmp: MINE1_EXPL_ROM_TYPE :=
  (
    "000000000000000110000000", --0
    "000000000000000110000000", --1
    "010000000100001110000000", --2
    "011100000110011110000000", --3
    "001110000111011110000000", --4
    "001111101111111111111000", --5
    "000111111111111111110000", --6
    "000011111111111111110000", --7
    "000111111111111111111111", --8
    "111111111111111111111111", --9
    "011111111111111111111100", --10
    "001111111111111111111000", --11
    "000111111111111111111100", --12
    "000111111111111111111111", --13
    "001111111111111111111111", --14
    "111111111111111111110000", --15
    "000000111111111111110000", --16
    "000000111111111101110000", --17
    "000001110111111100110000", --18
    "000001100111011100011000", --19
    "000000000110001100000000", --20
    "000000000110001100000000", --21
    "000000000110000000000000", --22
    "000000000100000000000000"  --23
  );
  signal mine10_expl_rom_addr: unsigned(4 downto 0);
  signal mine10_expl_rom_col: unsigned(4 downto 0);
  signal mine10_expl_rom_data: std_logic_vector(23 downto 0);
  signal mine10_expl_rom_bit: std_logic;

  -- mine2 explosion
  type MINE2_EXPL_ROM_TYPE is array (0 to 31) of std_logic_vector(31 downto 0);
  constant mine20_expl_bmp: MINE2_EXPL_ROM_TYPE :=
  (
    "00000000000000000000010000000000", --0
    "00000000000000000000110000000000", --1
    "00000000000000000000110000000000", --2
    "01000000000011000001110000000000", --3
    "01110000000011000011110000000000", --4
    "00111100000011100011110000000000", --5
    "00011111000111110111110001110000", --6
    "00001111100111111111111111110000", --7
    "00001111111111111111111111100000", --8
    "00000111111111111111111111000000", --9
    "00000011111111111111111111000000", --10
    "00001111111111111111111111111111", --11
    "11111111111111111111111111111111", --12
    "01111111111111111111111111111100", --13
    "00111111111111111111111111111000", --14
    "00011111111111111111111111100000", --15
    "00001111111111111111111111111000", --16
    "00000111111111111111111111111100", --17
    "00001111111111111111111111111111", --18
    "00111111111111111111111111111111", --19
    "01111111111111111111111111000000", --20
    "01110000111111111111111111000000", --21
    "00000000111111111111101111100000", --22
    "00000000111111111111100111100000", --23
    "00000001111011110111100011100000", --24
    "00000001100011100111100001100000", --25
    "00000000000011100011100000100000", --26
    "00000000000011100011100000000000", --27
    "00000000000011100001100000000000", --28
    "00000000000011000000000000000000", --29
    "00000000000011000000000000000000", --30
    "00000000000011000000000000000000"  --31
  );
  signal mine20_expl_rom_addr: unsigned(4 downto 0);
  signal mine20_expl_rom_col: unsigned(4 downto 0);
  signal mine20_expl_rom_data: std_logic_vector(31 downto 0);
  signal mine20_expl_rom_bit: std_logic;
  
 
  -- Tunnel Object
  type STATE_TYPE_TUNNEL is (NEW_GAME, PLAY, GAME_OVER_MESSAGE);
  signal state_tunnel_reg, state_tunnel_next: STATE_TYPE_TUNNEL;
  signal graphics_still: std_logic := '1'; -- freeze everything during new game or game over
  constant TUNNEL_WIDTH : integer:=1280;
  constant TUNNEL_HEIGHT : integer:=480; 
  constant TUNNEL_DELTA_V: integer:=1; -- speed of moving "camera" to the right over tunnel bmp
  signal actual_tunnel_on: std_logic; 
  -- tunnel_bmp
  signal tunnel_addr_row: unsigned(8 downto 0); -- need 9 bits to index 480 rows
  signal tunnel_addr_column: unsigned (10 downto 0); -- need 11 bits to index 1280 columns
  signal tunnel_bit: std_logic;
  -- tunnel "moving window" left and right tile indices;
  -- wraps around the tunnel_bmp;
  signal tunnel_l_reg, tunnel_l_next : unsigned(10 downto 0);
  signal tunnel_r_reg, tunnel_r_next : unsigned(10 downto 0);
  
  
begin

  -- (pixel_x,pixel_y) scan constantly the frame of 640x480; our job here is
  -- to see what we should display at that location - by checking 
  -- if coordinates are inside the ship area, tunnel, missile, mines, etc.
  pix_x <= unsigned(pixel_x);
  pix_y <= unsigned(pixel_y);
  
  
  -- registers Ship, Missile, Mines
  process (clk, reset, graphics_still)
  begin
    if (reset='1' or graphics_still='1') then -- graphics_still keeps all as if reset is applied to bring mines off the screen
      ship_x_reg <= (OTHERS=>'0');
      ship_y_reg <= to_unsigned((MAX_Y-SHIP_HEIGHT)/2,10); -- place Ship in the middle of screen on y axis;
      missile_x_reg <= (OTHERS=>'0'); 
      missile_y_reg <= (OTHERS=>'0');
      mine10_x_reg <= to_unsigned(MAX_X,10); -- right edge of screen horizontally
      mine10_y_reg <= to_unsigned((MAX_Y-MINE1_HEIGHT)/2,10); -- middle of screen vertically
      mine20_x_reg <= to_unsigned(MAX_X,10); -- right edge of screen horizontally
      mine20_y_reg <= to_unsigned((MAX_Y-MINE2_HEIGHT)/2,10); -- middle of screen vertically
    elsif (clk'event and clk='1') then
      ship_x_reg <= ship_x_next;
      ship_y_reg <= ship_y_next;     
      missile_x_reg <= missile_x_next;
      missile_y_reg <= missile_y_next;
      mine10_x_reg <= mine10_x_next;
      mine10_y_reg <= mine10_y_next;
      mine20_x_reg <= mine20_x_next;
      mine20_y_reg <= mine20_y_next;
    end if;
  end process;
  

  --===========================================================================================================================
  -- TUNNEL 
  
  -- instantiate countdown timer
  -- we use it to insert a delay of 4 sec to show the game over message;
  timer_4sec_in_tunnel_U0: entity work.timer
    generic map(W=>7) -- 4 seconds timer
    port map(clk=>clk, reset=>reset,
            timer_tick=>countdown_timer_tick,
            timer_start=>timer_4sec_start,
            timer_up=>timer_4sec_up);  


  -- Tunnel object main FSM
  -- (1) registers
  process (clk, reset) -- 50 MHz
  begin
    if reset='1' then
       state_tunnel_reg <= NEW_GAME;
    elsif (clk'event and clk='1') then
       state_tunnel_reg <= state_tunnel_next;
    end if;
  end process;
  
  -- (2) next-state logic
  process(game_over_from_ship, btn, timer_4sec_up, state_tunnel_reg) 
  begin
    state_tunnel_next <= state_tunnel_reg;  
    in_state_new_game <= '0';
    in_state_game_over_message <= '0';
    graphics_still <= '1'; -- freeze graphics
    timer_4sec_start <='0';    
    case state_tunnel_reg is
      when NEW_GAME =>
        in_state_new_game <= '1';
        if (btn(1)='1' or btn(0)='1') then -- buttons up/down pressed means player wants to start a new game 
          state_tunnel_next <= PLAY;
        end if;
      when PLAY =>
        graphics_still <= '0'; -- animated screen
        if (game_over_from_ship='1') then
          state_tunnel_next <= GAME_OVER_MESSAGE;
          timer_4sec_start <= '1'; -- 4 sec timer
        end if;
      when GAME_OVER_MESSAGE =>
        in_state_game_over_message <= '1';
        -- wait for 4 sec to display game over
        if timer_4sec_up='1' then
          state_tunnel_next <= NEW_GAME;
        end if;
      end case;
  end process;
  
  
  -- we use a moving window or "camera" that is 480x680 pixels and moving to the right
  -- with wrapping around when it gets to the right hand side of tunnel_bmp
  -- (1) registers 
  process (TIME_TICK, reset, graphics_still)
  begin
    if (reset='1' or graphics_still='1') then
      tunnel_l_reg <= "00000000000"; --0
      tunnel_r_reg <= "00111011111"; --479
      missile_x0_explosion_reg <= (OTHERS=>'0');
      ship_x0_explosion_reg <= (OTHERS=>'0');
      mine10_x0_explosion_reg <= (OTHERS=>'0');
      mine20_x0_explosion_reg <= (OTHERS=>'0');
    elsif (TIME_TICK'event and TIME_TICK='1') then
      tunnel_l_reg <= tunnel_l_next;
      tunnel_r_reg <= tunnel_r_next;
      missile_x0_explosion_reg <= missile_x0_explosion_next;
      ship_x0_explosion_reg <= ship_x0_explosion_next;
      mine10_x0_explosion_reg <= mine10_x0_explosion_next;
      mine20_x0_explosion_reg <= mine20_x0_explosion_next;
    end if;
  end process;
  
  -- (2) logic
  process (tunnel_l_reg, tunnel_r_reg, graphics_still,
    ship_x0_explosion_reg, 
    missile_x0_explosion_reg,
    mine10_x0_explosion_reg, mine20_x0_explosion_reg)
  begin 
    -- track ship location all the time; when hits wall, freeze it on Tunnel  
    ship_x0_explosion_next <= ship_x_reg; 
    if (explode_ship='1') then
      ship_x0_explosion_next <= ship_x0_explosion_reg - TUNNEL_DELTA_V; 
    end if;   
    -- track missile location all the time; when hits wall OR hits mine20 1st time only
    -- we freeze it on Tunnel, so that it "moves" together with Tunnel to left;
    missile_x0_explosion_next <= missile_x_reg; 
    if (explode_missile='1') then
      missile_x0_explosion_next <= missile_x0_explosion_reg - TUNNEL_DELTA_V; 
    end if;
    -- track mine10 location all the time; when it is hit by missile or ship, freeze it on Tunnel
    -- for explosion purposes
    mine10_x0_explosion_next <= mine10_x_reg; 
    if (explode_mine10='1') then
      mine10_x0_explosion_next <= mine10_x0_explosion_reg - TUNNEL_DELTA_V; 
    end if;
    -- track mine20 location all the time; when it is hit by missile or ship, freeze it on Tunnel
    -- for explosion purposes
    mine20_x0_explosion_next <= mine20_x_reg; 
    if (explode_mine20='1') then
      mine20_x0_explosion_next <= mine20_x0_explosion_reg - TUNNEL_DELTA_V; 
    end if;
    
    if (tunnel_l_reg < TUNNEL_WIDTH) then
      tunnel_l_next <= tunnel_l_reg + 1;
    else
      tunnel_l_next <= (OTHERS=>'0');
    end if;
    if (tunnel_r_reg < TUNNEL_WIDTH) then
      tunnel_r_next <= tunnel_r_reg + 1;
    else
      tunnel_r_next <= (OTHERS=>'0');
    end if; 
    if (graphics_still='1') then -- new game situation, hold still till user triggers
      tunnel_l_next <= "00000000000"; --0
      tunnel_r_next <= "00111011111"; --479
    end if;
  end process;  
  

  -- the Tunnel moving-window is always on screen, but, only the 
  -- top and bottom parts really are tunnel walls, rest is empty space;
  tunnel_addr_row    <= pix_y(8 downto 0); 
  tunnel_addr_column <= 
    (tunnel_l_reg + unsigned('0'&pix_x(9 downto 0))) when (tunnel_l_reg + unsigned('0'&pix_x(9 downto 0)))<TUNNEL_WIDTH else
    (tunnel_l_reg + unsigned('0'&pix_x(9 downto 0))) - TUNNEL_WIDTH; 
  
  -- instantiate Tunnel ROM
  tunnel_walls_unit: entity work.tunnel_rom
    port map(
      addr_row => tunnel_addr_row,
      addr_column => tunnel_addr_column, 
      tunnel_bit => tunnel_bit 
    );
  actual_tunnel_on <= '1' when (tunnel_bit='1') else '0';
  tunnel_rgb <= "100"; -- red



  --===========================================================================================================================
  -- SHIP object 
  
  TIME_TICK <= vsync; -- Ship takes as clock the TIME_TICK, 1/30 sec
  
  take_off_ev <= '1' when (btn(2)='1' or btn(1)='1' or btn(0)='1') else '0'; -- user starts Game; NOT really used
  player_ship_move <= '1' when (btn(1)='1' or btn(0)='1') else '0'; -- user moves ship down or up?
  player_fire_missile <= btn(2); -- essentially fire Missile, will be passed as fire_missile to Missile object
  
  ship_hit_mine <= ship_hit_mine_from_mine10 or ship_hit_mine_from_mine20; -- ship hit a mine: mine10 OR mine20, event sent to Ship object;
  
  
  ship_unit: entity work.ship
    port map(
      reset=> (reset or graphics_still),
      clk=>clk, -- 50 MHz clock
      countdown_timer_tick=>countdown_timer_tick,
      TIME_TICK=>TIME_TICK, -- clock of 30 cycles per second
      btn=>btn, -- pass to Ship also the actual button controls
      PLAYER_FIRE => player_fire_missile,
      PLAYER_SHIP_MOVE => player_ship_move, -- event that comes with coordinates info
      TAKE_OFF => take_off_ev, -- event generated by Tunnel when Player starts game
      score_val => score_total_val, -- score value passed with event SCORE 
      SCORE => score_ev, -- event generated
      x => ship_curr_x, -- passed with event SHIP_IMG
      y => ship_curr_y, -- passed with event SHIP_IMG
      ship_flying=> ship_is_flying, -- true when ship is flying
      SHIP_IMG => ship_img_ev, -- event posted to Tunnel
      HIT_MINE => ship_hit_mine, -- event posted by Tunnel from Mine1 or Mine2; Ship will explode
      mine_type => mine_type_hit, -- actually we have just 2 types of mines
      HIT_WALL => ship_hit_wall_ev_recorded, -- event posted by Tunnel; Ship will explode
      MISSILE_FIRE => fire_missile, -- event posted to Missile; includes x,y too
      DESTROYED_MINE => destroyed_mine_ev, -- event from Missile
      score_inc_val => score_delta_val_from_missile, -- how much to add to ship total score when mine is destroyed
      EXPLOSION_SHIP => explode_ship, -- event posted to Tunnel
      ship_explosion_size => ship_explosion_size, -- passed with event EXPLOSION_SHIP
      GAME_OVER => game_over_from_ship
    );     
  -- is current pixel inside the square bounding box of ship? 
  ship_x_l <= ship_x_reg;
  ship_y_t <= ship_y_reg;
  ship_x_r <= ship_x_l + SHIP_WIDTH - 1;
  ship_y_b <= ship_y_t + SHIP_HEIGHT - 1;
  bbox_ship_on <=
    '1' when (ship_x_l<=pix_x) and (pix_x<=ship_x_r) and
             (ship_y_t<=pix_y) and (pix_y<=ship_y_b) else
    '0';
  -- once inside the rectangular bbox of ship, is pixel actually ship pixel or background? 
  ship_rom_addr <= (pix_y(4 downto 0) - ship_y_t(4 downto 0)) when (bbox_ship_on='1') else "00000";
  ship_rom_col  <= (pix_x(5 downto 0) - ship_x_l(5 downto 0)) when (bbox_ship_on='1') else "000000";
  ship_rom_data <= ship_bmp(to_integer(ship_rom_addr));
  ship_rom_bit  <= ship_rom_data(SHIP_WIDTH-1 - to_integer(ship_rom_col));
  actual_ship_on <=
    '1' when (bbox_ship_on='1') and (ship_rom_bit='1') else
    '0';
  ship_rgb <= "100"; -- red
  -- new Ship position
  ship_y_next <= unsigned(ship_curr_y); 
  ship_x_next <= 
    (unsigned(ship_curr_x))           when (explode_ship='0') else 
    (unsigned(ship_x0_explosion_reg)) when (explode_ship='1') else 
    ship_x_reg;   
  
  
  --===========================================================================================================================  
  -- MISSILE object 

  missile_hit_mine <= missile_hit_mine10_ev_recorded or missile_hit_mine20_ev_recorded; -- missile hit a mine: mine10 OR mine20, event recorded is sent to Missile object; 
  
  missile_destroyed_mine <= missile_destroyed_mine10 or missile_destroyed_mine20; -- missile destroyed a mine: mine10 OR mine20, event sent to Missile object; 
  score_delta_destroyed_mine_1_or_2 <=  -- passed to Missile object, which will pass to Ship object
    std_logic_vector(to_unsigned(SCORE_DELTA_FOR_MINE1,20)) when (missile_destroyed_mine10='1') else -- 20
    std_logic_vector(to_unsigned(SCORE_DELTA_FOR_MINE2,20)) when (missile_destroyed_mine20='1') else -- 50
    (OTHERS=>'0');

  
  missile_unit: entity work.missile
    port map(
      reset=>(reset or graphics_still), -- reset or graphics_still or game_over_from_ship
      clk=>clk, -- 50 MHz clock
      countdown_timer_tick=>countdown_timer_tick,
      TIME_TICK=>TIME_TICK, -- clock of 30 cycles per second
      MISSILE_FIRE=> fire_missile, -- btn(2)
      x0 => std_logic_vector(ship_x_reg + MISSILE_WIDTH), -- pass ship x location to Missile object
      y0 => std_logic_vector(ship_y_reg), -- pass ship y location to Missile object
      x => missile_curr_x, -- passed with event MISSILE_IMG
      y => missile_curr_y, -- passed with event MISSILE_IMG
      missile_flying=> missile_is_flying, -- true when missile in flight
      DESTROYED_EITHER_MINE=> missile_destroyed_mine, -- event posted by Tunnel
      HIT_MINE=> missile_hit_mine, -- event posted by Tunnel to Missile object
      score_from_mine=> score_delta_destroyed_mine_1_or_2, -- score value from Tunnel to Missile object, with event HIT_MINE   
      HIT_MINE2_1ST_TIME=> missile_hit_mine20_1st_time, -- event from mine20 to missile via Tunnel
      HIT_WALL=> missile_hit_wall_ev_recorded, -- event posted by Tunnel
      MISSILE_IMG=> missile_IMG_ev, -- event posted to Tunnel; includes x,y too
      DESTROYED_MINE=> destroyed_mine_ev, -- event posted to Ship
      score_val=> score_delta_val_from_missile, -- score value passed with event SCORE to Ship (essentially what comes from Mines, via Missile, sent to Ship)
      EXPLOSION_MISSILE=> explode_missile, -- event posted to Tunnel
      missile_explosion_size=> missile_explosion_size -- passed with event EXPLOSION_MISSILE    
    );

  -- is current pixel inside the square bounding box of missile?
  missile_x_l <= missile_x_reg;
  missile_y_t <= missile_y_reg;
  missile_x_r <= missile_x_l + MISSILE_WIDTH - 1;
  missile_y_b <= missile_y_t + MISSILE_HEIGHT - 1;
  bbox_missile_on <=
    '1' when (missile_x_l<=pix_x) and (pix_x<=missile_x_r) and
             (missile_y_t<=pix_y) and (pix_y<=missile_y_b) else
    '0';
  -- once inside the rectangular bbox of missile, is pixel actually Missile pixel or background? 
  missile_rom_addr <= (pix_y(2 downto 0) - missile_y_t(2 downto 0)) when (bbox_missile_on='1') else "000";
  missile_rom_col  <= (pix_x(3 downto 0) - missile_x_l(3 downto 0)) when (bbox_missile_on='1') else "0000";
  missile_rom_data <= missile_bmp(to_integer(missile_rom_addr));
  missile_rom_bit <= missile_rom_data(MISSILE_WIDTH-1 - to_integer(missile_rom_col)); 
  actual_missile_on <=
    '1' when (bbox_missile_on='1') and (missile_rom_bit='1') and (missile_is_flying='1') else
    '0';
  missile_rgb <= "100"; -- red
  -- missile position; get it from the Missile object, which internally does the updates;
  -- missile moves horizontally till hitting something or out of screen area;
  missile_y_next <= (unsigned(missile_curr_y)+SHIP_HEIGHT-MISSILE_HEIGHT) when missile_is_flying='1' else 
    missile_y_reg;
  missile_x_next <= 
    (unsigned(missile_curr_x))           when (missile_is_flying='1' and explode_missile='0') else 
    (unsigned(missile_x0_explosion_reg)) when (missile_is_flying='0' and explode_missile='1') else 
    missile_x_reg;  

   

  --===========================================================================================================================  
  -- MINES objects 
  
  game_exit_from_user <= '0';
  
  -- --------------------------------------------------------------------------------------------------------------------------
  -- -----------------------------------------------Type 1 Mine Objects 
  -- mine10, mine11, mine12, ... for now we use only one mine of type 1
  
  recycle_mine10 <= '0';

  mine10: entity work.mine1 
    generic map(ID=> 0)
    port map(
      reset=>(reset or graphics_still), -- reset or graphics_still or game_over_from_ship
      clk=>clk, -- 50 MHz clock
      countdown_timer_tick=>countdown_timer_tick,
      TIME_TICK=>TIME_TICK, -- clock of 30 cycles per second NOT -- clk_10Hz,
      x0 => std_logic_vector(mine10_x_rand), -- pass random mine10 x location to Mine object
      y0 => std_logic_vector(mine10_y_rand), 
      MINE1_PLANT=>plant_mine10,
      MINE1_RECYCLE=>recycle_mine10,
      MINE1_IMG=>mine10_is_planted, -- event generated to Tunnel
      mine1_bmp_overlaps_ship_bmp=> ship_hit_mine10_ev_recorded, -- from checker of collision recorder of Ship with Mine1; tell Mine object; will take it and pass it tot Ship
      HIT_MINE1=> ship_hit_mine_from_mine10, -- event generated to Ship via Tunnel, will cause Ship to explode, mine to dissapear
      mine1_bmp_overlaps_missile_bmp=> missile_hit_mine10_ev_recorded, -- from checker of collision recorder of Missile with Mine1 object
      DESTROYED_MINE1=> missile_destroyed_mine10, -- event generated to Missile
      EXPLOSION_MINE1=> explode_mine10, -- event generated to Tunnel
      exit_action=> game_exit_from_user, -- from Player
      MINE1_DISABLED=> mine10_disabled, -- event generated to Tunnel
      mine1_id=> mine10_id, -- info passed with event MINE1_DISABLED
      x => mine10_curr_x, -- passed with event MISSILE_IMG
      y => mine10_curr_y, -- passed with event MISSILE_IMG
      mine1_explosion_size=> mine10_explosion_size
    );  
  
  -- is current pixel inside the square bounding box of mine10?
  mine10_x_l <= mine10_x_reg;
  mine10_y_t <= mine10_y_reg;
  mine10_x_r <= mine10_x_l + MINE1_WIDTH - 1;
  mine10_y_b <= mine10_y_t + MINE1_HEIGHT - 1;
  bbox_mine10_on <=
    '1' when (mine10_is_planted='1') and 
             (mine10_x_l<=pix_x) and (pix_x<=mine10_x_r) and
             (mine10_y_t<=pix_y) and (pix_y<=mine10_y_b) else
    '0';
  -- once inside the rectangular bbox of mine10, is pixel actually mine10 pixel or background? 
  mine10_rom_addr <= (pix_y(4 downto 0) - mine10_y_t(4 downto 0)) when (bbox_mine10_on='1') else "00000";
  mine10_rom_col  <= (pix_x(4 downto 0) - mine10_x_l(4 downto 0)) when (bbox_mine10_on='1') else "00000";
  mine10_rom_data <= mine10_bmp(to_integer(mine10_rom_addr));
  mine10_rom_bit <= mine10_rom_data(MINE1_WIDTH-1 - to_integer(mine10_rom_col)); 
  actual_mine10_on <=
    '1' when (bbox_mine10_on='1') and (mine10_rom_bit='1') else
    '0';
  mine10_rgb <= "011";
  -- mine10 moves horizontally to left, at the speed of Tunnel, because
  -- inside the tunnel the mine is fixed; it moves to left to create
  -- the illusion of ship moving to right; 
  -- it moves to left until it is destroyed, or hits the ship, or left wall and gets out
  -- mine10 position: get it from the Mine1 object, which internally does the updates upto an explosion;
  mine10_y_next <= (unsigned(mine10_curr_y)) when mine10_is_planted='1' else 
    mine10_y_reg;
  mine10_x_next <= 
    (unsigned(mine10_curr_x))           when (mine10_is_planted='1' and explode_mine10='0') else 
    (unsigned(mine10_x0_explosion_reg)) when (mine10_is_planted='0' and explode_mine10='1') else 
    mine10_x_reg;

  -- am I looking at a pixel inside area around mine10 with 32 pixels larger
  -- in all directions? I do not want to place mine20 in this area, to avoid mines overlap!
  bbox_expanded_mine10_on <=
    '1' when (mine10_is_planted='1') and 
             (mine10_x_l<=(pix_x+32)) and (pix_x<=(mine10_x_r+32)) and
             (mine10_y_t<=(pix_y+32)) and (pix_y<=(mine10_y_b+32)) else
    '0';
    
  
  -- --------------------------------------------------------------------------------------------------------------------------
  -- -----------------------------------------------Type 2 Mine Objects
  -- mine20, mine21, mine22, ... for now we use only one mine of type 2
  
  recycle_mine20 <= '0';

  mine20: entity work.mine2 
    generic map(ID=> 0)
    port map(
      reset=>(reset or graphics_still), -- reset or graphics_still or game_over_from_ship
      clk=>clk, -- 50 MHz clock
      countdown_timer_tick=>countdown_timer_tick,
      TIME_TICK=>TIME_TICK, -- clock of 30 cycles per second NOT -- clk_10Hz,
      x0 => std_logic_vector(mine20_x_rand), -- pass random mine20 x location to Mine object
      y0 => std_logic_vector(mine20_y_rand), 
      MINE2_PLANT=>plant_mine20,
      MINE2_RECYCLE=>recycle_mine20,
      MINE2_IMG=>mine20_is_planted, -- event generated to Tunnel
      mine2_bmp_overlaps_ship_bmp=> ship_hit_mine20_ev_recorded, -- from checker of collision recorder of Ship with Mine2; tell Mine object; will take it and pass it tot Ship
      HIT_MINE2=> ship_hit_mine_from_mine20, -- event generated to Ship via Tunnel, will cause Ship to explode, mine to dissapear
      mine2_bmp_overlaps_missile_bmp=> missile_hit_mine20_ev_recorded, -- from checker of collision recorder of Missile with Mine2 object
      mine2_hit_1st_time=> missile_hit_mine20_1st_time, -- event generated by mine2 for missile, passed via Tunnel
      DESTROYED_MINE2=> missile_destroyed_mine20, -- event generated to Missile
      EXPLOSION_MINE2=> explode_mine20, -- event generated to Tunnel     
      exit_action=> game_exit_from_user, -- from Player
      MINE2_DISABLED=> mine20_disabled, -- event generated to Tunnel
      mine2_id=> mine20_id, -- info passed with event MINE2_DISABLED
      x => mine20_curr_x, -- passed with event MISSILE_IMG
      y => mine20_curr_y, -- passed with event MISSILE_IMG
      mine2_explosion_size=> mine20_explosion_size
    );  
  
  -- is current pixel inside the square bounding box of mine20?
  mine20_x_l <= mine20_x_reg;
  mine20_y_t <= mine20_y_reg;
  mine20_x_r <= mine20_x_l + MINE2_WIDTH - 1;
  mine20_y_b <= mine20_y_t + MINE2_HEIGHT - 1;
  bbox_mine20_on <=
    '1' when (mine20_is_planted='1') and 
             (mine20_x_l<=pix_x) and (pix_x<=mine20_x_r) and
             (mine20_y_t<=pix_y) and (pix_y<=mine20_y_b) else
    '0';
  -- once inside the rectangular bbox of mine20, is pixel actually mine20 pixel or background? 
  mine20_rom_addr <= (pix_y(4 downto 0) - mine20_y_t(4 downto 0)) when (bbox_mine20_on='1') else "00000";
  mine20_rom_col  <= (pix_x(4 downto 0) - mine20_x_l(4 downto 0)) when (bbox_mine20_on='1') else "00000";
  mine20_rom_data <= mine20_bmp(to_integer(mine20_rom_addr));
  mine20_rom_bit <= mine20_rom_data(MINE2_WIDTH-1 - to_integer(mine20_rom_col)); 
  actual_mine20_on <=
    '1' when (bbox_mine20_on='1') and (mine20_rom_bit='1') else
    '0';
  mine20_rgb <= "010";
  -- mine20 moves horizontally to left, at the speed of Tunnel, because
  -- inside the tunnel the mine is fixed; it moves to left to create
  -- the illusion of ship moving to right; 
  -- it moves to left until it is destroyed, or hits the ship, or left wall and gets out
  -- mine20 position: get it from the Mine1 object, which internally does the updates upto an explosion;
  mine20_y_next <= (unsigned(mine20_curr_y)) when mine20_is_planted='1' else 
    mine20_y_reg;
  mine20_x_next <= 
    (unsigned(mine20_curr_x))           when (mine20_is_planted='1' and explode_mine20='0') else 
    (unsigned(mine20_x0_explosion_reg)) when (mine20_is_planted='0' and explode_mine20='1') else 
    mine20_x_reg;
  
  -- am I looking at a pixel inside area around mine20 with 24 pixels larger
  -- in all directions? I do not want to place mine10 in this area, to avoid mines overlap!
  bbox_expanded_mine20_on <=
    '1' when (mine20_is_planted='1') and
             (mine20_x_l<=(pix_x+24)) and (pix_x<=(mine20_x_r+24)) and
             (mine20_y_t<=(pix_y+24)) and (pix_y<=(mine20_y_b+24)) else
    '0';
    

  -- --------------------------------------------------------------------------------------------------------------------------
  -- -----------------------------------------------logic to plant mines
  
  -- use LFSRs to generate lots of pseudorandom numbers, 0-1024;
  -- use those as potential locations to place mines;
  
  -- instantiate countdown timer
  -- used to provide random seed to the first LFSR; sampled at time
  -- user presses button "Up"; in this way we insert "user-randomness" into the
  -- "pseudorandomness" of the LFSR; 
  counter_rollover_U0: entity work.counter_rollover
    port map(clk=>clk, reset=>reset, sample_now=>btn(0), z=>seed_for_LFSR);
            
  -- instantiate 4 LFSRs on 10 bits, 2 for mine10 locations and 2 for mine20 locations
  -- for mine10 locations
  inst_lfsr10_mine10_x: entity work.lfsr10
    port map(
      reset=>reset, -- reset or graphics_still or game_over_from_ship
      clk=>TIME_TICK, -- NOTE: during a TIME_TICK, we scan all pixels on screen! during scanning I will have once (x_rand=pix_x and y_rand=pix_y)
      seed => seed_for_LFSR, -- different for any different run of the game!
      z => x_rand_lfsr_mine10 -- random x location; 
    ); 
  inst_lfsr10_mine10_y: entity work.lfsr10 
    port map(
      reset=>reset, 
      clk=>TIME_TICK, 
      seed => "1111111111",
      z => y_rand_lfsr_mine10 -- random y location;
    ); 
  -- for mine20 locations
  inst_lfsr10_mine20_x: entity work.lfsr10
    port map(
      reset=>reset, 
      clk=>pixel_tick, 
      seed => "0000011111",
      z => x_rand_lfsr_mine20  
    ); 
  inst_lfsr10_mine20_y: entity work.lfsr10 
    port map(
      reset=>reset, 
      clk=>pixel_tick,
      seed => "1100110011",
      z => y_rand_lfsr_mine20 
    ); 
    
  -- 1) out of those random numbers, we should pick up only qualifyable locations to plant mines;
  -- locations should not be on wall areas, and should not be placed too close to Ship
  -- use a band guard of 200 pixels; also, mines should not overlap;
  process (pixel_tick, reset, graphics_still) -- clk
  begin
    if (reset='1') then --or graphics_still='1'
      mine10_x_rand_reg <= to_unsigned((MAX_X-MINE1_WIDTH)/2,10); -- place mine10 in the middle of screen on x axis;
      mine10_y_rand_reg <= to_unsigned((MAX_Y-MINE1_HEIGHT)/2,10); -- place mine10 in the middle of screen on y axis;
      mine20_x_rand_reg <= to_unsigned(MAX_X,10); -- place mine20 on the right edge of screen on x axis;
      mine20_y_rand_reg <= to_unsigned((MAX_Y-MINE2_HEIGHT)/2,10); -- place mine10 in the middle of screen on y axis;  
    elsif (pixel_tick'event and pixel_tick='1') then
      mine10_x_rand_reg <= mine10_x_rand_next; 
      mine10_y_rand_reg <= mine10_y_rand_next;   
      mine20_x_rand_reg <= mine20_x_rand_next; 
      mine20_y_rand_reg <= mine20_y_rand_next;
    end if;
  end process; 
  -- 2) logic to always record and keep available valid locations
  -- to plant mines; this good locations generator provide locations 
  -- for both types of mines;  
  process (
    pix_x, pix_y,
    x_rand_lfsr_mine10, y_rand_lfsr_mine10, 
    x_rand_lfsr_mine20, y_rand_lfsr_mine20,
    actual_tunnel_on, 
    bbox_expanded_mine10_on, bbox_expanded_mine20_on,
    mine10_x_rand_reg, mine10_y_rand_reg, 
    mine20_x_rand_reg, mine20_y_rand_reg)
  begin 
    mine10_x_rand_next <= mine10_x_rand_reg; 
    mine10_y_rand_next <= mine10_y_rand_reg;
    mine20_x_rand_next <= mine20_x_rand_reg; 
    mine20_y_rand_next <= mine20_y_rand_reg;    
    -- NOTE: during a TIME_TICK, we scan all pixels on screen! during scanning I will have for sure 
    -- once: (x_rand=pix_x and y_rand=pix_y); when this happens and the location is not good,
    -- we look the next random location and so on; each new random loc is generated at 1/30 sec rate
    -- withing one such interval, all pixels are scanned
    if (x_rand_lfsr_mine10=pix_x and y_rand_lfsr_mine10=pix_y) then
      if (actual_tunnel_on='0' and bbox_expanded_mine20_on='0' and x_rand_lfsr_mine10>128) then -- not on wall or in vicity of mine20; to right of a band
        mine10_x_rand_next <= x_rand_lfsr_mine10;
        mine10_y_rand_next <= y_rand_lfsr_mine10;
      end if;
    end if;
    
    if (x_rand_lfsr_mine20=pix_x and y_rand_lfsr_mine20=pix_y) then
      if (actual_tunnel_on='0' and bbox_expanded_mine10_on='0' and x_rand_lfsr_mine20>256) then -- not on wall or in vicity of mine10; to right of a band
        mine20_x_rand_next <= x_rand_lfsr_mine20;
        mine20_y_rand_next <= y_rand_lfsr_mine20;
      end if;
    end if;
  end process;
  
  

  -- logic to plant mines
  process (TIME_TICK, reset)
  begin
    if (reset = '1') then 
      plant_mine_state_reg <= PLANT_PAUSE;
    elsif (TIME_TICK' event and TIME_TICK = '1') then 
      plant_mine_state_reg <= plant_mine_state_next;
    end if;
  end process; 
  
  process (plant_mine_state_reg,
    mine10_x_rand_reg, mine10_y_rand_reg,
    mine20_x_rand_reg, mine20_y_rand_reg)
  begin 
    plant_mine_state_next <= plant_mine_state_reg;
    plant_mine10 <= '0';
    plant_mine20 <= '0';
    
    case plant_mine_state_reg is 
      when PLANT_PAUSE =>
        plant_mine_state_next <= PLANT_MINE1;
      when PLANT_MINE1 =>
        if (mine10_is_planted='0') then
          mine10_x_rand <= mine10_x_rand_reg;
          mine10_y_rand <= mine10_y_rand_reg;
          plant_mine10 <= '1';
          plant_mine_state_next <= PLANT_MINE2;
        end if;
      when PLANT_MINE2 =>
        if (mine20_is_planted='0') then
          mine20_x_rand <= mine20_x_rand_reg;
          mine20_y_rand <= mine20_y_rand_reg;
          plant_mine20 <= '1';
          plant_mine_state_next <= PLANT_MINE1;
        end if;
    end case;
  end process;   
  

  --===========================================================================================================================  
  -- COLLISION DETECTION logic
  ship_hit_wall_ev <= 
    '1' when (actual_ship_on='1' and actual_tunnel_on='1') else 
    '0';
  ship_hit_mine10_ev <= 
    '1' when (actual_ship_on='1' and actual_mine10_on='1') else 
    '0'; 
  ship_hit_mine20_ev <= 
    '1' when (actual_ship_on='1' and actual_mine20_on='1') else 
    '0'; 
  missile_hit_wall_ev <= 
    '1' when (actual_missile_on='1' and actual_tunnel_on='1') else 
    '0';
  missile_hit_mine10_ev <= 
    '1' when (actual_missile_on='1' and actual_mine10_on='1') else 
    '0';
  missile_hit_mine20_ev <= 
    '1' when (actual_missile_on='1' and actual_mine20_on='1') else 
    '0';    
    
  -- Events sent to Ship must be synchronized with TIME_TICK clock - the clock
  -- that all UML statechrts use to operate; the pixels sweeping happens at clk frequncy,
  -- much higher; difference in this timing may make pixel-overlap-events (used
  -- to detect collisions) to go unnoticed; they may be too short and not be "seen" by 
  -- the UML inside Ship; that is why these collision "recorders" records a collison 
  -- situation and keeps it till the next clock edge of the TIME_TICK "clock signal" for Ship object;
  collision_ship_tunnel_unit: entity work.collision_recorder
    port map(
      clk=>clk, reset=>reset,
      clear=>TIME_TICK, -- we want at the end of frame to know all collisions 
      pixels_overlap_event=>ship_hit_wall_ev,
      collision_detected=>ship_hit_wall_ev_recorded);   

  -- recorder of collision between Ship and mine10
  collision_ship_mine10_unit: entity work.collision_recorder
    port map(
      clk=>clk, reset=>reset,
      clear=>TIME_TICK, -- we want at the end of frame to know all collisions 
      pixels_overlap_event=>ship_hit_mine10_ev,
      collision_detected=>ship_hit_mine10_ev_recorded);  

  -- recorder of collision between Ship and mine20
  collision_ship_mine20_unit: entity work.collision_recorder
    port map(
      clk=>clk, reset=>reset,
      clear=>TIME_TICK, -- we want at the end of frame to know all collisions 
      pixels_overlap_event=>ship_hit_mine20_ev,
      collision_detected=>ship_hit_mine20_ev_recorded); 
      
  -- recorder of collision between missile and wall
  collision_missile_tunnel_unit: entity work.collision_recorder
    port map(
      clk=>clk, reset=>reset,
      clear=>TIME_TICK, -- we want at the end of frame to know all collisions 
      pixels_overlap_event=>missile_hit_wall_ev,
      collision_detected=>missile_hit_wall_ev_recorded);
      
  -- recorder of collision between missile and mine10
  collision_missile_mine10_unit: entity work.collision_recorder
    port map(
      clk=>clk, reset=>reset,
      clear=>TIME_TICK, -- we want at the end of frame to know all collisions 
      pixels_overlap_event=>missile_hit_mine10_ev,
      collision_detected=>missile_hit_mine10_ev_recorded); 

  -- recorder of collision between missile and mine20
  collision_missile_mine20_unit: entity work.collision_recorder
    port map(
      clk=>clk, reset=>reset,
      clear=>TIME_TICK, -- we want at the end of frame to know all collisions 
      pixels_overlap_event=>missile_hit_mine20_ev,
      collision_detected=>missile_hit_mine20_ev_recorded);  


  --===========================================================================================================================
  -- EXPLOSIONS 
  
  -- Ship explodes when hits wall
  -- once inside the rectangular bbox of ship, is pixel actually ship-explosion pixel or background? 
  ship_expl_rom_addr <= (pix_y(4 downto 0) - ship_y_t(4 downto 0)) when (bbox_ship_on='1') else "00000";
  ship_expl_rom_col  <= (pix_x(5 downto 0) - ship_x_l(5 downto 0)) when (bbox_ship_on='1') else "000000";
  ship_expl_rom_data <= ship_expl_bmp(to_integer(ship_rom_addr));
  ship_expl_rom_bit  <= ship_expl_rom_data(SHIP_WIDTH-1 - to_integer(ship_expl_rom_col));
  actual_ship_expl_on <=
    '1' when (bbox_ship_on='1') and (ship_expl_rom_bit='1') else
    '0';
  ship_expl_rgb <= "001"; -- blue
  
  
  -- Missile, when hits wall
  -- is current pixel inside the square bounding box of missile-explossion?
  -- NOTE: I make the explosion to be larger than the missile itself
  -- missile is 8x16 and the explosion is 8 pixels larger in all directions: 24x32
  missile_expl_x_l <= missile_x_reg - 8;
  missile_expl_y_t <= missile_y_reg - 8;
  missile_expl_x_r <= missile_expl_x_l + MISSILE_EXPL_WIDTH - 1;
  missile_expl_y_b <= missile_expl_y_t + MISSILE_EXPL_HEIGHT - 1;
  bbox_missile_expl_on <=
    '1' when (missile_expl_x_l<=pix_x) and (pix_x<=missile_expl_x_r) and
             (missile_expl_y_t<=pix_y) and (pix_y<=missile_expl_y_b) else
    '0';
  -- once inside the rectangular bbox of missile explosion, is pixel actually Missile Explosion pixel or background? 
  missile_expl_rom_addr <= (pix_y(4 downto 0) - missile_expl_y_t(4 downto 0)) when (bbox_missile_expl_on='1') else "00000";
  missile_expl_rom_col  <= (pix_x(4 downto 0) - missile_expl_x_l(4 downto 0)) when (bbox_missile_expl_on='1') else "00000";
  missile_expl_rom_data <= missile_expl_bmp(to_integer(missile_expl_rom_addr));
  missile_expl_rom_bit <= missile_expl_rom_data(MISSILE_EXPL_WIDTH-1 - to_integer(missile_expl_rom_col)); 
  actual_missile_expl_on <=
    '1' when (bbox_missile_expl_on='1') and (missile_expl_rom_bit='1')  else 
    '0';
  missile_expl_rgb <= "001"; -- blue  
  
  
  -- Mine1, when is hit by Missile
  -- is current pixel inside the square bounding box of mine10 explosion bbox?
  mine10_expl_x_l <= mine10_x_reg;
  mine10_expl_y_t <= mine10_y_reg;
  mine10_expl_x_r <= mine10_expl_x_l + MINE1_WIDTH - 1;
  mine10_expl_y_b <= mine10_expl_y_t + MINE1_HEIGHT - 1;
  bbox_expl_mine10_on <=
    '1' when (mine10_expl_x_l<=pix_x) and (pix_x<=mine10_expl_x_r) and
             (mine10_expl_y_t<=pix_y) and (pix_y<=mine10_expl_y_b) else
    '0';
  -- once inside the rectangular bbox of mine10 explosion, is pixel actually Mine1 Explosion pixel or background? 
  mine10_expl_rom_addr <= (pix_y(4 downto 0) - mine10_y_t(4 downto 0)) when (bbox_expl_mine10_on='1') else "00000";
  mine10_expl_rom_col  <= (pix_x(4 downto 0) - mine10_x_l(4 downto 0)) when (bbox_expl_mine10_on='1') else "00000";
  mine10_expl_rom_data <= mine10_expl_bmp(to_integer(mine10_expl_rom_addr));
  mine10_expl_rom_bit <= mine10_expl_rom_data(MINE1_WIDTH-1 - to_integer(mine10_expl_rom_col)); 
  actual_mine10_expl_on <=
    '1' when (bbox_expl_mine10_on='1') and (mine10_expl_rom_bit='1')  else 
    '0';
  mine10_expl_rgb <= "001"; -- blue  
 
 
  -- Mine2, when is hit by Missile - TWICE!
  -- is current pixel inside the square bounding box of mine20 explosion bbox?
  mine20_expl_x_l <= mine20_x_reg;
  mine20_expl_y_t <= mine20_y_reg;
  mine20_expl_x_r <= mine20_expl_x_l + MINE2_WIDTH - 1;
  mine20_expl_y_b <= mine20_expl_y_t + MINE2_HEIGHT - 1;
  bbox_expl_mine20_on <=
    '1' when (mine20_expl_x_l<=pix_x) and (pix_x<=mine20_expl_x_r) and
             (mine20_expl_y_t<=pix_y) and (pix_y<=mine20_expl_y_b) else
    '0';
  -- once inside the rectangular bbox of mine20 explosion, is pixel actually Mine1 Explosion pixel or background? 
  mine20_expl_rom_addr <= (pix_y(4 downto 0) - mine20_y_t(4 downto 0)) when (bbox_expl_mine20_on='1') else "00000";
  mine20_expl_rom_col  <= (pix_x(4 downto 0) - mine20_x_l(4 downto 0)) when (bbox_expl_mine20_on='1') else "00000";
  mine20_expl_rom_data <= mine20_expl_bmp(to_integer(mine20_expl_rom_addr));
  mine20_expl_rom_bit <= mine20_expl_rom_data(MINE2_WIDTH-1 - to_integer(mine20_expl_rom_col)); 
  actual_mine20_expl_on <=
    '1' when (bbox_expl_mine20_on='1') and (mine20_expl_rom_bit='1')  else 
    '0';
  mine20_expl_rgb <= "001"; -- blue   
  
  
  --===========================================================================================================================  
  -- rgb multiplexing circuit
  process(
    explode_ship,
    actual_tunnel_on,   
    bbox_mine10_on, actual_mine10_on, bbox_expl_mine10_on, actual_mine10_expl_on,
    bbox_mine20_on, actual_mine20_on, bbox_expl_mine20_on, actual_mine20_expl_on,
    actual_missile_on, bbox_missile_expl_on, actual_missile_expl_on,
    bbox_ship_on, actual_ship_on, actual_ship_expl_on,
    tunnel_rgb, 
    mine10_rgb, mine10_expl_rgb,
    mine20_rgb, mine20_expl_rgb,
    missile_rgb, missile_expl_rgb,
    ship_rgb, ship_expl_rgb) 
  begin
    rgb <= "110"; -- yellow background

    if (actual_tunnel_on='1') then     
      rgb <= tunnel_rgb;
    end if;    

    if (bbox_mine10_on='1' or bbox_expl_mine10_on='1') then
      if (explode_mine10='1') then
        if (actual_mine10_expl_on='1') then
          rgb <= mine10_expl_rgb;
        end if;
      else -- mine10 is not exploding
        if (actual_mine10_on='1') then
          rgb <= mine10_rgb;
        end if;
      end if;
    end if;    

    if (bbox_mine20_on='1'  or bbox_expl_mine20_on='1') then
      if (explode_mine20='1') then
        if (actual_mine20_expl_on='1') then
          rgb <= mine20_expl_rgb;
        end if;
      else -- mine20 is not exploding
        if (actual_mine20_on='1') then
          rgb <= mine20_rgb;
        end if;
      end if;
    end if;
    
    if (actual_missile_on='1') then    
      rgb <= missile_rgb;
    end if;    
    if (bbox_missile_expl_on='1') then
      if (explode_missile='1') then
        if (actual_missile_expl_on='1') then
          rgb <= missile_expl_rgb;
        end if;
      end if;
    end if;
    
    if (bbox_ship_on='1') then
      if (explode_ship='1') then
        if (actual_ship_expl_on='1') then
          rgb <= ship_expl_rgb;
        end if;
      else -- ship is not exploding
        if (actual_ship_on='1') then
          rgb <= ship_rgb;
        end if;
      end if;
    end if;
 
  end process;

  -- graphics on display? update graph_on signal
  graph_on <= 
    actual_tunnel_on or 
    actual_mine10_on or actual_mine10_expl_on or
    actual_mine20_on or actual_mine20_expl_on or
    actual_ship_on or actual_ship_expl_on or 
    actual_missile_on or actual_missile_expl_on; 
    
  -- overall score so far;
  score <= score_total_val; -- score_total_val comes from Ship object; passed here to out port to top level, which will pass it to game_text
  
end arch;