library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity ship is
  port(
    reset: in std_logic; 
    clk: in std_logic; -- 50 MHz clock; used for count-down timers only
    countdown_timer_tick: in std_logic; -- used by 2 sec and 4 sec countdown timers
    TIME_TICK: in std_logic; -- clock of 30 cycles per second; main clock for Ship
    btn: std_logic_vector(2 downto 0); -- KEY2: fire Missile; KEY1,0: Ship down/up;
    PLAYER_FIRE: in std_logic; -- player fires missile
    PLAYER_SHIP_MOVE: in std_logic; -- event that comes with coordinates info
    TAKE_OFF: in std_logic; -- event generated by Tunnel when Player starts game
    score_val: out std_logic_vector(19 downto 0); -- score value passed with event SCORE 
    SCORE: out std_logic; -- event generated
    x, y: out std_logic_vector(9 downto 0); -- passed with event SHIP_IMG
    ship_flying: out std_logic; -- true when ship is flying
    SHIP_IMG: out std_logic; -- event posted to Tunnel
    HIT_MINE: in std_logic; -- event posted by Tunnel 
    mine_type: in std_logic_vector(1 downto 0); -- actually we have just 2 types of mines
    HIT_WALL: in std_logic; -- event posted by Tunnel
    MISSILE_FIRE: out std_logic; -- event posted to Missile; includes x,y too
    DESTROYED_MINE: in std_logic; -- event from Missile
    score_inc_val: in std_logic_vector(19 downto 0); -- how much to add to local score when mine is destroyed
    EXPLOSION_SHIP: out std_logic; -- event posted to Tunnel
    ship_explosion_size: out std_logic_vector(9 downto 0); -- passed with event EXPLOSION_SHIP
    GAME_OVER: out std_logic
  );
end ship;


architecture UML_ARCHITECTURE of ship is

  type SUPERSTATE_TYPE_SHIP is (ACTIVE, INACTIVE);
  type STATE_TYPE_SHIP is (Parked, Flying, Exploding);
  signal superstate_reg, superstate_next : SUPERSTATE_TYPE_SHIP;
  signal state_reg, state_next : STATE_TYPE_SHIP;
  -- coordinates 
  signal x_reg, x_next: unsigned(9 downto 0);
  signal y_reg, y_next: unsigned(9 downto 0); 
  signal score_reg, score_next: unsigned(19 downto 0);
  signal local_ctr_reg, local_ctr_next: unsigned(7 downto 0); -- local counter; count TIME_TICK 30 times (i.e., 1 sec) and increment score
  signal exp_ctr_reg, exp_ctr_next: unsigned(9 downto 0); -- explosion counter
  signal timer_2sec_start, timer_2sec_up: std_logic;
  
  constant MAX_X: integer:=640;
  constant MAX_Y: integer:=480;
  constant SHIP_HEIGHT : integer:=32;
  constant SHIP_DELTA_V: integer:=2; -- displacement to move on move-upp or move-down
  
  begin
  
    -- state register; process #1
    process (TIME_TICK, reset)
    begin
      if (reset = '1') then 
        superstate_reg <= INACTIVE;
        state_reg <= Parked;
        x_reg <= (OTHERS=>'0');
        y_reg <= to_unsigned((MAX_Y-SHIP_HEIGHT)/2,10); -- place Ship in the middle of screen on y axis;
        score_reg <= (OTHERS=>'0');
        local_ctr_reg <= (OTHERS=>'0');
      elsif (TIME_TICK' event and TIME_TICK = '1') then 
        superstate_reg <= superstate_next;
        state_reg <= state_next;
        x_reg <= x_next;
        y_reg <= y_next;
        score_reg <= score_next;
        local_ctr_reg <= local_ctr_next;
      end if;
    end process;   
    
    -- next state and output logic; process #2
    process (superstate_reg, state_reg, exp_ctr_reg, 
      PLAYER_FIRE, PLAYER_SHIP_MOVE, TAKE_OFF, 
      DESTROYED_MINE, HIT_MINE, HIT_WALL)
    begin
      -- default initializations
      superstate_next <= superstate_reg;
      state_next <= state_reg;
      x_next <= x_reg;
      y_next <= y_reg;
      score_next <= score_reg;
      local_ctr_next <= local_ctr_reg;
      ship_flying<='0'; 
      SCORE <= '0';
      SHIP_IMG <= '0';
      MISSILE_FIRE <= '0';
      EXPLOSION_SHIP <= '0';
      GAME_OVER <= '0';
      timer_2sec_start <='0';     

      case superstate_reg is 
        --=====================================================================
        when INACTIVE => -- superstate
          --if PLAYER_FIRE = '1' then
          
          if PLAYER_SHIP_MOVE = '1' then
            superstate_next <= ACTIVE;
            --x_next <= unsigned(x0);
            --y_next <= unsigned(y0);
          end if; 
        --=====================================================================
        when ACTIVE => -- superstate; all action happens here! 
          case state_reg is 
            --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
            when Parked =>
              -- place Ship at default, initial location
              x_next <= (OTHERS=>'0'); 
              y_next <= to_unsigned((MAX_Y-SHIP_HEIGHT)/2,10);
              if PLAYER_SHIP_MOVE = '1' then -- Player starts game
                state_next <= Flying;
                score_next <= (OTHERS=>'0'); -- reset score
                SCORE <= '1'; -- generate event SCORE upon entry into Flying state
                local_ctr_next <= (OTHERS=>'0'); -- reset local counter (counts 0-9)
              end if;
            --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
            when Flying => 
              if btn(1)='1' and (y_reg + SHIP_HEIGHT - 1)<(MAX_Y-1-SHIP_DELTA_V) then
                y_next <= y_reg + SHIP_DELTA_V; -- move down
              elsif btn(0)='1' and y_reg>SHIP_DELTA_V then
                y_next <= y_reg - SHIP_DELTA_V; -- move up
              end if;
              
              ship_flying<='1';
              SHIP_IMG <= '1'; -- generate event SHIP_IMG; passed with coordinates info
              local_ctr_next <= local_ctr_reg + 1; 
              if (local_ctr_reg = 30)  then
                score_next <= score_reg + 1; -- increment score for surviving another second in the game
                SCORE <= '1'; -- generate event SCORE to Tunnel to update score
                local_ctr_next <= (OTHERS=>'0'); -- reset local counter
              end if;
              if PLAYER_FIRE = '1' then
                MISSILE_FIRE <= '1'; -- generate event MISSILE_FIRE to Missile object
              end if;
              if DESTROYED_MINE = '1' then
                -- add to local score the amount passed thru event; amount which depends
                -- on the type of mine destroyed;
                score_next <= score_reg + unsigned(score_inc_val); 
              end if;
              if (HIT_MINE = '1' or HIT_WALL = '1') then
                state_next <= Exploding;
                exp_ctr_next <= (OTHERS=>'0'); -- clear explosion counter
                timer_2sec_start <='1'; -- start cowntdown counter 2 sec
              end if;
            --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~                
            when Exploding =>  
              EXPLOSION_SHIP <= '1'; -- post event to Tunnel
              -- wait for 2 sec to display exploding ship
              if timer_2sec_up='1' then
                state_next <= Parked;
                GAME_OVER <= '1'; -- generate event to Tunnel
                superstate_next <= INACTIVE; 
              end if;             
            --~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
          end case; 
        --=====================================================================  
      end case;
    end process;
 
  -- score passed with event SCORE generated by Ship
  score_val <= std_logic_vector(score_reg);
  
  -- coordinates passed with events SHIP_IMG
  x <= std_logic_vector(x_reg);
  y <= std_logic_vector(y_reg); 
  
  -- instantiate countdown timer
  timer_2sec_U0: entity work.timer
    generic map(W=>6) -- 2 seconds timer
    port map(clk=>clk, reset=>reset,
            timer_tick=>countdown_timer_tick,
            timer_start=>timer_2sec_start,
            timer_up=>timer_2sec_up);
  
end UML_ARCHITECTURE;  
